// float_1.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module float_1 (
		input  wire        s1_clk,    // s1.clk
		input  wire        s1_clk_en, //   .clk_en
		input  wire [31:0] s1_dataa,  //   .dataa
		input  wire [31:0] s1_datab,  //   .datab
		input  wire [1:0]  s1_n,      //   .n
		input  wire        s1_reset,  //   .reset
		input  wire        s1_start,  //   .start
		output wire        s1_done,   //   .done
		output wire [31:0] s1_result  //   .result
	);

	fpoint_wrapper #(
		.useDivider (0)
	) nios_custom_instr_floating_point_0 (
		.clk    (s1_clk),    // s1.clk
		.clk_en (s1_clk_en), //   .clk_en
		.dataa  (s1_dataa),  //   .dataa
		.datab  (s1_datab),  //   .datab
		.n      (s1_n),      //   .n
		.reset  (s1_reset),  //   .reset
		.start  (s1_start),  //   .start
		.done   (s1_done),   //   .done
		.result (s1_result)  //   .result
	);

endmodule
