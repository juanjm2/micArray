// Audio_config.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module Audio_config (
		input  wire  audio_and_video_config_0_clk_clk,                 //                audio_and_video_config_0_clk.clk
		inout  wire  audio_and_video_config_0_external_interface_SDAT, // audio_and_video_config_0_external_interface.SDAT
		output wire  audio_and_video_config_0_external_interface_SCLK, //                                            .SCLK
		input  wire  audio_and_video_config_0_reset_reset              //              audio_and_video_config_0_reset.reset
	);

	Audio_config_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (audio_and_video_config_0_clk_clk),                 //                    clk.clk
		.reset       (audio_and_video_config_0_reset_reset),             //                  reset.reset
		.address     (),                                                 // avalon_av_config_slave.address
		.byteenable  (),                                                 //                       .byteenable
		.read        (),                                                 //                       .read
		.write       (),                                                 //                       .write
		.writedata   (),                                                 //                       .writedata
		.readdata    (),                                                 //                       .readdata
		.waitrequest (),                                                 //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT), //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)  //                       .export
	);

endmodule
