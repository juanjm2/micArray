module fifo_play(
	input logic sck,
	input logic record,
	input logic play,
	input logic [31:0] left_channel,
	input logic [31:0] right_channel,
);

endmodule
