// float.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module float (
		input  wire        clk_clk,                                           //                                     clk.clk
		input  wire [31:0] nios_custom_instr_floating_point_2_0_s1_dataa,     // nios_custom_instr_floating_point_2_0_s1.dataa
		input  wire [31:0] nios_custom_instr_floating_point_2_0_s1_datab,     //                                        .datab
		input  wire [3:0]  nios_custom_instr_floating_point_2_0_s1_n,         //                                        .n
		output wire [31:0] nios_custom_instr_floating_point_2_0_s1_result,    //                                        .result
		input  wire        nios_custom_instr_floating_point_2_0_s2_clk,       // nios_custom_instr_floating_point_2_0_s2.clk
		input  wire        nios_custom_instr_floating_point_2_0_s2_clk_en,    //                                        .clk_en
		input  wire [31:0] nios_custom_instr_floating_point_2_0_s2_dataa,     //                                        .dataa
		input  wire [31:0] nios_custom_instr_floating_point_2_0_s2_datab,     //                                        .datab
		input  wire [2:0]  nios_custom_instr_floating_point_2_0_s2_n,         //                                        .n
		input  wire        nios_custom_instr_floating_point_2_0_s2_reset,     //                                        .reset
		input  wire        nios_custom_instr_floating_point_2_0_s2_reset_req, //                                        .reset_req
		input  wire        nios_custom_instr_floating_point_2_0_s2_start,     //                                        .start
		output wire        nios_custom_instr_floating_point_2_0_s2_done,      //                                        .done
		output wire [31:0] nios_custom_instr_floating_point_2_0_s2_result,    //                                        .result
		input  wire        reset_reset_n                                      //                                   reset.reset_n
	);

	float_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (nios_custom_instr_floating_point_2_0_s1_dataa),     // s1.dataa
		.s1_datab     (nios_custom_instr_floating_point_2_0_s1_datab),     //   .datab
		.s1_n         (nios_custom_instr_floating_point_2_0_s1_n),         //   .n
		.s1_result    (nios_custom_instr_floating_point_2_0_s1_result),    //   .result
		.s2_clk       (nios_custom_instr_floating_point_2_0_s2_clk),       // s2.clk
		.s2_clk_en    (nios_custom_instr_floating_point_2_0_s2_clk_en),    //   .clk_en
		.s2_dataa     (nios_custom_instr_floating_point_2_0_s2_dataa),     //   .dataa
		.s2_datab     (nios_custom_instr_floating_point_2_0_s2_datab),     //   .datab
		.s2_n         (nios_custom_instr_floating_point_2_0_s2_n),         //   .n
		.s2_reset     (nios_custom_instr_floating_point_2_0_s2_reset),     //   .reset
		.s2_reset_req (nios_custom_instr_floating_point_2_0_s2_reset_req), //   .reset_req
		.s2_start     (nios_custom_instr_floating_point_2_0_s2_start),     //   .start
		.s2_done      (nios_custom_instr_floating_point_2_0_s2_done),      //   .done
		.s2_result    (nios_custom_instr_floating_point_2_0_s2_result)     //   .result
	);

endmodule
