module gain(
);

endmodule
