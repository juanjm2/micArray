
module Audio_config (
	audio_and_video_config_0_clk_clk,
	audio_and_video_config_0_reset_reset,
	audio_and_video_config_0_external_interface_SDAT,
	audio_and_video_config_0_external_interface_SCLK);	

	input		audio_and_video_config_0_clk_clk;
	input		audio_and_video_config_0_reset_reset;
	inout		audio_and_video_config_0_external_interface_SDAT;
	output		audio_and_video_config_0_external_interface_SCLK;
endmodule
