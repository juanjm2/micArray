
module audio_pll (
	audio_pll_0_audio_clk_clk,
	audio_pll_0_ref_clk_clk,
	audio_pll_0_ref_reset_reset,
	audio_pll_0_reset_source_reset);	

	output		audio_pll_0_audio_clk_clk;
	input		audio_pll_0_ref_clk_clk;
	input		audio_pll_0_ref_reset_reset;
	output		audio_pll_0_reset_source_reset;
endmodule
