// aud_24.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module aud_24 (
		input  wire        clk_clk,                //              clk.clk
		input  wire        ext_ADCDAT,             //              ext.ADCDAT
		input  wire        ext_ADCLRCK,            //                 .ADCLRCK
		input  wire        ext_BCLK,               //                 .BCLK
		output wire        ext_DACDAT,             //                 .DACDAT
		input  wire        ext_DACLRCK,            //                 .DACLRCK
		inout  wire        ext_1_SDAT,             //            ext_1.SDAT
		output wire        ext_1_SCLK,             //                 .SCLK
		input  wire [15:0] fir_left_input_data,    //   fir_left_input.data
		input  wire        fir_left_input_valid,   //                 .valid
		input  wire [1:0]  fir_left_input_error,   //                 .error
		output wire [23:0] fir_left_output_data,   //  fir_left_output.data
		output wire        fir_left_output_valid,  //                 .valid
		output wire [1:0]  fir_left_output_error,  //                 .error
		input  wire [15:0] fir_right_input_data,   //  fir_right_input.data
		input  wire        fir_right_input_valid,  //                 .valid
		input  wire [1:0]  fir_right_input_error,  //                 .error
		output wire [23:0] fir_right_output_data,  // fir_right_output.data
		output wire        fir_right_output_valid, //                 .valid
		output wire [1:0]  fir_right_output_error, //                 .error
		input  wire [23:0] left_input_data,        //       left_input.data
		input  wire        left_input_valid,       //                 .valid
		output wire        left_input_ready,       //                 .ready
		input  wire        left_output_ready,      //      left_output.ready
		output wire [23:0] left_output_data,       //                 .data
		output wire        left_output_valid,      //                 .valid
		input  wire        reset_reset_n,          //            reset.reset_n
		input  wire [23:0] right_input_data,       //      right_input.data
		input  wire        right_input_valid,      //                 .valid
		output wire        right_input_ready,      //                 .ready
		input  wire        right_output_ready,     //     right_output.ready
		output wire [23:0] right_output_data,      //                 .data
		output wire        right_output_valid      //                 .valid
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [FIR_LEFT:reset_n, FIR_RIGHT:reset_n, audio_0:reset, audio_and_video_config_0:reset]

	aud_24_FIR_LEFT fir_left (
		.clk              (clk_clk),                         //                     clk.clk
		.reset_n          (~rst_controller_reset_out_reset), //                     rst.reset_n
		.ast_sink_data    (fir_left_input_data),             //   avalon_streaming_sink.data
		.ast_sink_valid   (fir_left_input_valid),            //                        .valid
		.ast_sink_error   (fir_left_input_error),            //                        .error
		.ast_source_data  (fir_left_output_data),            // avalon_streaming_source.data
		.ast_source_valid (fir_left_output_valid),           //                        .valid
		.ast_source_error (fir_left_output_error)            //                        .error
	);

	aud_24_FIR_LEFT fir_right (
		.clk              (clk_clk),                         //                     clk.clk
		.reset_n          (~rst_controller_reset_out_reset), //                     rst.reset_n
		.ast_sink_data    (fir_right_input_data),            //   avalon_streaming_sink.data
		.ast_sink_valid   (fir_right_input_valid),           //                        .valid
		.ast_sink_error   (fir_right_input_error),           //                        .error
		.ast_source_data  (fir_right_output_data),           // avalon_streaming_source.data
		.ast_source_valid (fir_right_output_valid),          //                        .valid
		.ast_source_error (fir_right_output_error)           //                        .error
	);

	aud_24_audio_0 audio_0 (
		.clk                          (clk_clk),                        //                         clk.clk
		.reset                        (rst_controller_reset_out_reset), //                       reset.reset
		.from_adc_left_channel_ready  (left_output_ready),              //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (left_output_data),               //                            .data
		.from_adc_left_channel_valid  (left_output_valid),              //                            .valid
		.from_adc_right_channel_ready (right_output_ready),             // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (right_output_data),              //                            .data
		.from_adc_right_channel_valid (right_output_valid),             //                            .valid
		.to_dac_left_channel_data     (left_input_data),                //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (left_input_valid),               //                            .valid
		.to_dac_left_channel_ready    (left_input_ready),               //                            .ready
		.to_dac_right_channel_data    (right_input_data),               //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (right_input_valid),              //                            .valid
		.to_dac_right_channel_ready   (right_input_ready),              //                            .ready
		.AUD_ADCDAT                   (ext_ADCDAT),                     //          external_interface.export
		.AUD_ADCLRCK                  (ext_ADCLRCK),                    //                            .export
		.AUD_BCLK                     (ext_BCLK),                       //                            .export
		.AUD_DACDAT                   (ext_DACDAT),                     //                            .export
		.AUD_DACLRCK                  (ext_DACLRCK)                     //                            .export
	);

	aud_24_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk_clk),                        //                    clk.clk
		.reset       (rst_controller_reset_out_reset), //                  reset.reset
		.address     (),                               // avalon_av_config_slave.address
		.byteenable  (),                               //                       .byteenable
		.read        (),                               //                       .read
		.write       (),                               //                       .write
		.writedata   (),                               //                       .writedata
		.readdata    (),                               //                       .readdata
		.waitrequest (),                               //                       .waitrequest
		.I2C_SDAT    (ext_1_SDAT),                     //     external_interface.export
		.I2C_SCLK    (ext_1_SCLK)                      //                       .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
