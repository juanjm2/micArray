// line_in.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module line_in (
		input  wire [23:0] audio_0_avalon_left_channel_sink_data,            //            audio_0_avalon_left_channel_sink.data
		input  wire        audio_0_avalon_left_channel_sink_valid,           //                                            .valid
		output wire        audio_0_avalon_left_channel_sink_ready,           //                                            .ready
		input  wire        audio_0_avalon_left_channel_source_ready,         //          audio_0_avalon_left_channel_source.ready
		output wire [23:0] audio_0_avalon_left_channel_source_data,          //                                            .data
		output wire        audio_0_avalon_left_channel_source_valid,         //                                            .valid
		input  wire [23:0] audio_0_avalon_right_channel_sink_data,           //           audio_0_avalon_right_channel_sink.data
		input  wire        audio_0_avalon_right_channel_sink_valid,          //                                            .valid
		output wire        audio_0_avalon_right_channel_sink_ready,          //                                            .ready
		input  wire        audio_0_avalon_right_channel_source_ready,        //         audio_0_avalon_right_channel_source.ready
		output wire [23:0] audio_0_avalon_right_channel_source_data,         //                                            .data
		output wire        audio_0_avalon_right_channel_source_valid,        //                                            .valid
		input  wire        audio_0_external_interface_ADCDAT,                //                  audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,               //                                            .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                  //                                            .BCLK
		output wire        audio_0_external_interface_DACDAT,                //                                            .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,               //                                            .DACLRCK
		inout  wire        audio_and_video_config_0_external_interface_SDAT, // audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK, //                                            .SCLK
		input  wire        clk_clk,                                          //                                         clk.clk
		input  wire        reset_reset_n                                     //                                       reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [audio_0:reset, audio_and_video_config_0:reset]

	line_in_audio_0 audio_0 (
		.clk                          (clk_clk),                                   //                         clk.clk
		.reset                        (rst_controller_reset_out_reset),            //                       reset.reset
		.from_adc_left_channel_ready  (audio_0_avalon_left_channel_source_ready),  //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (audio_0_avalon_left_channel_source_data),   //                            .data
		.from_adc_left_channel_valid  (audio_0_avalon_left_channel_source_valid),  //                            .valid
		.from_adc_right_channel_ready (audio_0_avalon_right_channel_source_ready), // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (audio_0_avalon_right_channel_source_data),  //                            .data
		.from_adc_right_channel_valid (audio_0_avalon_right_channel_source_valid), //                            .valid
		.to_dac_left_channel_data     (audio_0_avalon_left_channel_sink_data),     //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (audio_0_avalon_left_channel_sink_valid),    //                            .valid
		.to_dac_left_channel_ready    (audio_0_avalon_left_channel_sink_ready),    //                            .ready
		.to_dac_right_channel_data    (audio_0_avalon_right_channel_sink_data),    //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (audio_0_avalon_right_channel_sink_valid),   //                            .valid
		.to_dac_right_channel_ready   (audio_0_avalon_right_channel_sink_ready),   //                            .ready
		.AUD_ADCDAT                   (audio_0_external_interface_ADCDAT),         //          external_interface.export
		.AUD_ADCLRCK                  (audio_0_external_interface_ADCLRCK),        //                            .export
		.AUD_BCLK                     (audio_0_external_interface_BCLK),           //                            .export
		.AUD_DACDAT                   (audio_0_external_interface_DACDAT),         //                            .export
		.AUD_DACLRCK                  (audio_0_external_interface_DACLRCK)         //                            .export
	);

	line_in_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk_clk),                                          //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                   //                  reset.reset
		.address     (),                                                 // avalon_av_config_slave.address
		.byteenable  (),                                                 //                       .byteenable
		.read        (),                                                 //                       .read
		.write       (),                                                 //                       .write
		.writedata   (),                                                 //                       .writedata
		.readdata    (),                                                 //                       .readdata
		.waitrequest (),                                                 //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT), //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)  //                       .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
